parameter M=16;
parameter N=24;
parameter LATENCY=26;
