module lut_ov5640_rgb565_480_272(
	input[9:0]             lut_index,   //Look-up table address
	output reg[31:0]       lut_data     //Device address (8bit I2C address), register address, register data
);




24'h3103_11
24'h3008_82
24'h3008_42
24'h3103_03
24'h3017_ff
24'h3018_ff
24'h3034_1a
24'h3037_13
24'h3108_01
24'h3630_36
24'h3631_0e
24'h3632_e2
24'h3633_12
24'h3621_e0
24'h3704_a0
24'h3703_5a
24'h3715_78
24'h3717_01
24'h370b_60
24'h3705_1a
24'h3905_02
24'h3906_10
24'h3901_0a
24'h3731_12
24'h3600_08
24'h3601_33
24'h302d_60
24'h3620_52
24'h371b_20
24'h471c_50
24'h3a13_43
24'h3a18_00
24'h3a19_f8
24'h3635_13
24'h3636_03
24'h3634_40
24'h3622_01
24'h3c01_34
24'h3c04_28
24'h3c05_98
24'h3c06_00
24'h3c07_08
24'h3c08_00
24'h3c09_1c
24'h3c0a_9c
24'h3c0b_40
24'h3810_00
24'h3811_10
24'h3812_00
24'h3708_64
24'h4001_02
24'h4005_1a
24'h3000_00
24'h3004_ff
24'h300e_58
24'h302e_00
24'h4300_60
24'h501f_01
24'h440e_00
24'h5000_a7
24'h3a0f_30
24'h3a10_28
24'h3a1b_30
24'h3a1e_26
24'h3a11_60
24'h3a1f_14
24'h5800_23
24'h5801_14
24'h5802_0f
24'h5803_0f
24'h5804_12
24'h5805_26
24'h5806_0c
24'h5807_08
24'h5808_05
24'h5809_05
24'h580a_08
24'h580b_0d
24'h580c_08
24'h580d_03
24'h580e_00
24'h580f_00
24'h5810_03
24'h5811_09
24'h5812_07
24'h5813_03
24'h5814_00
24'h5815_01
24'h5816_03
24'h5817_08
24'h5818_0d
24'h5819_08
24'h581a_05
24'h581b_06
24'h581c_08
24'h581d_0e
24'h581e_29
24'h581f_17
24'h5820_11
24'h5821_11
24'h5822_15
24'h5823_28
24'h5824_46
24'h5825_26
24'h5826_08
24'h5827_26
24'h5828_64
24'h5829_26
24'h582a_24
24'h582b_22
24'h582c_24
24'h582d_24
24'h582e_06
24'h582f_22
24'h5830_40
24'h5831_42
24'h5832_24
24'h5833_26
24'h5834_24
24'h5835_22
24'h5836_22
24'h5837_26
24'h5838_44
24'h5839_24
24'h583a_26
24'h583b_28
24'h583c_42
24'h583d_ce
24'h5180_ff
24'h5181_f2
24'h5182_00
24'h5183_14
24'h5184_25
24'h5185_24
24'h5186_09
24'h5187_09
24'h5188_09
24'h5189_75
24'h518a_54
24'h518b_e0
24'h518c_b2
24'h518d_42
24'h518e_3d
24'h518f_56
24'h5190_46
24'h5191_f8
24'h5192_04
24'h5193_70
24'h5194_f0
24'h5195_f0
24'h5196_03
24'h5197_01
24'h5198_04
24'h5199_12
24'h519a_04
24'h519b_00
24'h519c_06
24'h519d_82
24'h519e_38
24'h5480_01
24'h5481_08
24'h5482_14
24'h5483_28
24'h5484_51
24'h5485_65
24'h5486_71
24'h5487_7d
24'h5488_87
24'h5489_91
24'h548a_9a
24'h548b_aa
24'h548c_b8
24'h548d_cd
24'h548e_dd
24'h548f_ea
24'h5490_1d
24'h5381_1e
24'h5382_5b
24'h5383_08
24'h5384_0a
24'h5385_7e
24'h5386_88
24'h5387_7c
24'h5388_6c
24'h5389_10
24'h538a_01
24'h538b_98
24'h5580_06
24'h5583_40
24'h5584_10
24'h5589_10
24'h558a_00
24'h558b_f8
24'h501d_40
24'h5300_08
24'h5301_30
24'h5302_10
24'h5303_00
24'h5304_08
24'h5305_30
24'h5306_08
24'h5307_16
24'h5309_08
24'h530a_30
24'h530b_04
24'h530c_06
24'h5025_00
24'h3008_02
24'h3035_11
24'h3036_8C
24'h3c07_08
_
_
_
_
_
24'h3820_41
24'h3821_01
_
24'h3820_42
24'h3821_01
_
24'h3820_43
24'h3821_01
_
24'h3820_40
24'h3821_01
_
_
24'h3814_31
24'h3815_31
24'h3800_00
24'h3801_00
24'h3802_00
24'h3803_04
24'h3804_0a
24'h3805_3f
24'h3806_07
24'h3807_9b
24'h3808_01
24'h3809_e0
24'h380a_01
24'h380b_10
24'h380c_07
24'h380d_68
24'h380e_03
24'h380f_d8
24'h3813_06
24'h3618_00
24'h3612_29
24'h3709_52
24'h370c_03
24'h3a02_17
24'h3a03_10
24'h3a14_17
24'h3a15_10
24'h4004_02
24'h3002_1c
24'h3006_c3
24'h4713_03
24'h4407_04
24'h460b_35
24'h460c_22
24'h4837_22
24'h3824_02
24'h5001_a3
24'h3503_00
24'h3016_02
24'h3b07_0a
24'h3b00_83
24'h3b00_00
24'hffff_ff
h0000,8'_h0


endmodule 